class Config;
  int nErrors;
endclass
