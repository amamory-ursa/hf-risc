typedef enum bit [6:0] {
  OPCD_LUI   = 7'b01_101_11,
  OPCD_AUIPC = 7'b00_101_11,
  OPCD_JAL   = 7'b11_011_11,
  OPCD_JALR  = 7'b11_001_11,
  BRANCH     = 7'b11_000_11,
  LOAD       = 7'b00_000_11,
  STORE      = 7'b01_000_11,
  OPP_IMM    = 7'b00_100_11,
  OP         = 7'b01_100_11,
  SYSTEM     = 7'b11_100_11
}  Opcode;

bit[31:0] OpcodeMask[Opcode];
initial begin
  OpcodeMask[OPCD_LUI]   = 32'b0000000_00000_00000_000_00000_1111111;
  OpcodeMask[OPCD_AUIPC] = 32'b0000000_00000_00000_000_00000_1111111;
  OpcodeMask[OPCD_JAL]   = 32'b0000000_00000_00000_000_00000_1111111;
  OpcodeMask[OPCD_JALR]  = 32'b0000000_00000_00000_111_00000_1111111;
  OpcodeMask[BRANCH]     = 32'b0000000_00000_00000_111_00000_1111111;
  OpcodeMask[LOAD]       = 32'b0000000_00000_00000_111_00000_1111111;
  OpcodeMask[STORE]      = 32'b0000000_00000_00000_111_00000_1111111;
  OpcodeMask[OPP_IMM]    = 32'b0000000_00000_00000_111_00000_1111111;
  OpcodeMask[OP]         = 32'b1111111_00000_00000_111_00000_1111111;
  OpcodeMask[SYSTEM]     = 32'b1111111_11111_11111_111_11111_1111111;
end

bit[31:0] OpcodeMask_SR_I
                      = 32'b1111111_00000_00000_111_00000_1111111;

typedef enum bit[31:0] {
  LUI    = 32'b0000000_00000_00000_000_00000_0110111,

  AUIPC  = 32'b0000000_00000_00000_000_00000_0010111,

  JAL    = 32'b0000000_00000_00000_000_00000_1101111,

  JALR   = 32'b0000000_00000_00000_000_00000_1100111,

  BEQ    = 32'b0000000_00000_00000_000_00000_1100011,
  BNE    = 32'b0000000_00000_00000_001_00000_1100011,
  BLT    = 32'b0000000_00000_00000_100_00000_1100011,
  BGE    = 32'b0000000_00000_00000_101_00000_1100011,
  BLTU   = 32'b0000000_00000_00000_110_00000_1100011,
  BGEU   = 32'b0000000_00000_00000_111_00000_1100011,

  LB     = 32'b0000000_00000_00000_000_00000_0000011,
  LH     = 32'b0000000_00000_00000_001_00000_0000011,
  LW     = 32'b0000000_00000_00000_010_00000_0000011,
  LBU    = 32'b0000000_00000_00000_100_00000_0000011,
  LHU    = 32'b0000000_00000_00000_101_00000_0000011,

  SB     = 32'b0000000_00000_00000_000_00000_0100011,
  SH     = 32'b0000000_00000_00000_001_00000_0100011,
  SW     = 32'b0000000_00000_00000_010_00000_0100011,

  ADDI   = 32'b0000000_00000_00000_000_00000_0010011,
  SLTI   = 32'b0000000_00000_00000_010_00000_0010011,
  SLTIU  = 32'b0000000_00000_00000_011_00000_0010011,
  XORI   = 32'b0000000_00000_00000_100_00000_0010011,
  ORI    = 32'b0000000_00000_00000_110_00000_0010011,
  ANDI   = 32'b0000000_00000_00000_111_00000_0010011,
  SLLI   = 32'b0000000_00000_00000_001_00000_0010011,
  SRLI   = 32'b0000000_00000_00000_101_00000_0010011,
  SRAI   = 32'b0100000_00000_00000_101_00000_0010011,

  ADD    = 32'b0000000_00000_00000_000_00000_0110011,
  SUB    = 32'b0100000_00000_00000_000_00000_0110011,
  SLL    = 32'b0000000_00000_00000_001_00000_0110011,
  SLT    = 32'b0000000_00000_00000_010_00000_0110011,
  SLTU   = 32'b0000000_00000_00000_011_00000_0110011,
  XOR    = 32'b0000000_00000_00000_100_00000_0110011,
  SRL    = 32'b0000000_00000_00000_101_00000_0110011,
  SRA    = 32'b0100000_00000_00000_101_00000_0110011,
  OR     = 32'b0000000_00000_00000_110_00000_0110011,
  AND    = 32'b0000000_00000_00000_111_00000_0110011,
  // FENCE = 32'b0000000_00000_00000_000_00000_0000000,
  // FENCE.I = 32'b0000000_00000_00000_000_00000_0000000,
  ECALL  = 32'b0000000_00000_00000_000_00000_1110011,
  EBREAK = 32'b0000001_00000_00000_000_00000_1110011
  // CSRRW = 32'b0000000_00000_00000_000_00000_0000000,
  // CSRRS = 32'b0000000_00000_00000_000_00000_0000000,
  // CSRRC = 32'b0000000_00000_00000_000_00000_0000000,
  // CSRRWI = 32'b0000000_00000_00000_000_00000_0000000,
  // CSRRSI = 32'b0000000_00000_00000_000_00000_0000000,
  // CSRRCI = 32'b0000000_00000_00000_000_00000_0000000,
} Instruction;
