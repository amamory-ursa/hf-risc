typedef struct {
  bit [31:0] [31:0] registers;
  bit [31:0] pc;
} Snapshot;
