module top;
	dummy_ag ag1();
	dummy_ag_IO ag2();
	scoreboard sb1();
	dummy_chk chk1();
endmodule

