module top;
	dummy_ag ag1();
	scoreboard sb1();
	dummy_chk chk1();
endmodule

